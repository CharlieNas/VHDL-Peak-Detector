-- TEAM B 