-- TEAM A